���Z     @  <   I�      �  &                                       
    0                                                    !   �   F� 	   ,          � Project@Options� -�   !�     7   \+ 	   -          � File@@Version2.1  � 1.1     (                                                          1   f   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access8                   .       ,       )       3       �      �T      �#      �7      ��     ߜ     �     �n     �n     ��     �     �     ''     (0     ))     *Y     +�     ,,     -�     .E     /�     0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �0    !� BuildAll!� 0!� Contents!� Copyright � ...!�  !�  !�@     � 1017   �  ��6W     �  �� Al   
  � Index�� P|"   �   D+�� 
� ( / H     � Topic@Index  �    �  	5   !�3 "Index", ( 511, 0, 511, 1023), , , (192,192,192), 0!�  $   , 0!�4 "Glossary", ( 0, 0, 511, 1023), , , (192,192,192), 0%   ,192,192), 0!�. "", ( 0, 511, 1023, 511), , , (192,192,192)&   ), , , (192,192,192), 0!�, "", ( 0, 0, 1023, 511), , , (192'    "Guana", , , , (192,192,192), 0!�- "", ( 64, 64, 832, 832(   r  �  	   -          � F1ProjectWindowsC-�  L !�    �  !�  !�  !�  !�  !�                                      *     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !+   �   �� 	   -          � F1ProjectButtonsZ -�   !�  �. #include "stdafx.h",Topic4, 0,<IDH_MainWindow>!�( �����,-     � 	   .          � F1ProjectGlossary� -�  	 !      !�                                                       /     !� 0!�  !�  !� 0!� 0!� No!�  !� Guana!� 1!�  !�  !�6    T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE              w  ��� �� ��� ����������� ������ ������ ����� � ���� ���, ��� 4   M'  �0 	   ,          � F1ProjectStyle2'-�  � !�OL    Title , MS Sans Serif ,  18 ,  120 ,  250 ,  40 ,  40 ,  1W  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�   ������� ����� ������;!�- /B /Just L /Text �������� �� �����8   1  t �� 
� + 2 K     � Topic@Contents  �    � 9    	  � 1000   �  ��9Z     �  �� Dr     � Contents:   �� S�     �  �� 	c(  �-�   !� /T N /Just M /Text Con;   tents!�C /L N /Jump Index /Link /Macro /Play /popup Main /Jd  ust L /Text Index!�P /L /Jump IDH_MainWindow /Link /Macro /   ����������������� ���� ����� ������������ ������, ���� ���>   elp\img\CUR_GU~1.BMP /Just L /Text ������������, � �������   ������� ������������ � ������� ������ �����.��������!�%/R     /Z N /Style /Just L!� /X /Style /Just L  
u �           ?        �  �� 	`�   N -�   !� /T N /Just L /Text Index!� �2   ��, ��� ��������� ����� �������, �� ������, ������ ��������Q   180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagrapB    60 ,  0 ,  0 ,  0 , None , !�J Paragraph , Arial ,  10 ,  C   , None , !�J Paragraph , Arial ,  10 ,  180 ,  250 ,  20 , D   aph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 E     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�J ParagrF    0 , -1 ,  0 , None , !�R Paragraph , MS Sans Serif ,  10 ,G   None , !�F Title , Arial ,  18 ,  120 ,  250 ,  40 ,  40 , H   e , Arial ,  18 ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , I    ,  120 ,  250 ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F TitlJ   ,  40 ,  40 ,  0 , -1 ,  0 , None , !�F Title , Arial ,  18K    , -1 ,  0 , Shade , !�F Title , Arial ,  18 ,  120 ,  250 N   ����, ������� ��� �����������. ������� ����������� ��������O   �� ������ �� ���������� ������, ������� ��� �����������. ��P    ������ ���������� � ������� �� ������ �������� �� ���������   �� ����� ��������� ������� "<<Jump to".!�% /H /Just M /Text�`   h , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , a    ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 , -1 ,  0 , None , !R     20 ,  0 , -1 , -1 , None , !�T Jump Label , MS Sans SerifS    None , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,T   ng , Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 ,U   80 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , None , !�L Sub HeadiV    ,  0 , -1 , -1 , None , !�L Sub Heading , Arial ,  12 ,  1W   e , !�L Sub Heading , Arial ,  12 ,  180 ,  250 ,  40 ,  20X    Arial ,  12 ,  180 ,  250 ,  40 ,  20 ,  0 , -1 , -1 , NonY     250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�L Sub Heading ,Z    ,  0 , -1 ,  0 , None , !�H Heading , Arial ,  12 ,  180 ,[    None , !�H Heading , Arial ,  12 ,  180 ,  250 ,  60 ,  20\   ng , Arial ,  12 ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 ,]   ,  180 ,  250 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�H Headi^   0 ,  20 ,  1 , -1 ,  0 , Shade , !�H Heading , Arial ,  12 _   None , !�Q Heading , MS Sans Serif ,  14 ,  180 ,  250 ,  6�p   �L Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10q   Footnote , Arial ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,b   ,  8 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H c   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial d   0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  180 ,  25e   N Mono Spaced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  f    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�g    20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spaced , Courierh   0 , None , !�N Mono Spaced , Courier ,  10 ,  180 ,  250 , i   ced , Courier ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  j   180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�N Mono Spak     10 ,  0 ,  0 , None , !�N Mono Spaced , Courier ,  10 ,  l    , !�L Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  20 ,m   rial ,  10 ,  180 ,  250 ,  20 ,  20 ,  10 ,  0 ,  0 , Nonen   250 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�L Jump Label , Ao    ,  0 ,  0 , None , !�L Jump Label , Arial ,  10 ,  180 ,  �     0 , None , !�H Footnote , Arial ,  8 ,  180 ,  250 ,  20 �    ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�r   ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , Arials    , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 t   Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Noneu     20 ,  60 ,  0 ,  0 ,  0 , None , !�R Bitmap Jump Label , v    None , !�R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,w   ph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 ,x    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap Paragray    ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 ,  180 , z   Paragraph , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0{    180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Q Bitmap |    0 ,  0 ,  0 , None , !�Q Bitmap Paragraph , Arial ,  10 , }   aragraph , MS Sans Serif ,  10 ,  180 ,  250 ,  20 ,  60 , ~   180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�Y Bitmap P   ,  60 ,  0 ,  0 ,  0 , None , !�H Footnote , Arial ,  8 ,  ��   R Bitmap Jump Label , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    0 , None , !�M Outline Node , Arial ,  10 ,  180 ,  250 , �   Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 , �    ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumerated �    0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 ,  180�   ated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R Enumer�    0 ,  0 ,  0 , None , !�R Enumerated Bullet , Arial ,  10 ,�   numerated Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 , �    10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�R E�   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet , Arial , �    0 ,  0 ,  0 , None , !�G Bullet , Arial ,  10 ,  180 ,  25�   one , !�G Bullet , Arial ,  10 ,  180 ,  250 ,  20 ,  60 , �    , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , N�     180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�G Bullet�    ,  0 ,  0 ,  0 , None , !�O Bullet , MS Sans Serif ,  10 ,��    10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Node , Arial �   ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  10 ,  180 ,  25�    , None , !�E Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   Line , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�     10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�E �   10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial ,�   0 , None , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  �    Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  �    440 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline�   0 ,  0 ,  0 ,  0 , None , !�M Outline Leaf , Arial ,  10 , �   e , !�M Outline Leaf , Arial ,  10 ,  440 ,  250 ,  10 ,  1�    Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�    250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M Outline Node ,�   ,  0 ,  0 , None , !�M Outline Node , Arial ,  10 ,  180 , �    Outline Node , Arial ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 �   ,  10 ,  180 ,  250 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�M��   0 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Line , Arial ,  1�   ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Arial ,  10 ,  18�    ,  0 , None , !�F Index , Arial ,  10 ,  180 ,  250 ,  20 �   !�F Index , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0�   al ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , �    ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Index , Ari�     60 ,  0 , -1 ,  0 , None , !�F Index , Arial ,  10 ,  180�    !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,�   ial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None ,�   0 ,  60 ,  0 , -1 ,  0 , None , !�S Index Letter Label , Ar�   e , !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,  2�    Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , Non�     20 ,  60 ,  0 , -1 ,  0 , None , !�S Index Letter Label ,�   None , !�S Index Letter Label , Arial ,  12 ,  180 ,  250 ,�   e , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , �   0 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�E Lin�   0 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�V Glossary L�   mage , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0�    10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F I�   ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary , Arial , �     0 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 ,  250 �   !�I Glossary , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,�   al ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , �    250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�I Glossary , Ari�     0 , -1 ,  0 , None , !�I Glossary , Arial ,  10 ,  180 , �   sary Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,�    ,  180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glos�    , -1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12�   y Letter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0�    180 ,  250 ,  20 ,  60 ,  0 , -1 ,  0 , None , !�V Glossar�   -1 ,  0 , None , !�V Glossary Letter Label , Arial ,  12 , �   etter Label , Arial ,  12 ,  180 ,  250 ,  20 ,  60 ,  0 , :�    , None , !�F Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60�    , !�F Table , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,�   Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None�   180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , �   0 ,  60 ,  0 ,  0 ,  0 , None , !�F Table , Arial ,  10 ,  �    0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 ,  2�   e , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 , �    Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , Non�   ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar ,�    ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 �   ,  0 ,  0 ,  0 , None , !�D Bar , Arial ,  10 ,  180 ,  250�   0 , None , !�D Bar , Arial ,  10 ,  180 ,  250 ,  20 ,  60 �   Image , Arial ,  10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  �     10 ,  180 ,  250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F �   250 ,  20 ,  60 ,  0 ,  0 ,  0 , None , !�F Image , Arial ,�    ,  0 ,  0 ,  0 , None , !�F Image , Arial ,  10 ,  180 ,  6�     0 ,  0 , None , !�F Table , Arial ,  10 ,  180 ,  250 ,  �   0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  �    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 , �     ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,�   Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1�   �1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , �   ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�    ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �    0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0�    0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 , �     0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,�    ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 �    0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0�   20 ,  60 ,  0 ,  0 ,  0 , None , !�;  , Arial ,  10 ,  0 , ��   0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 �   ����� ��� ������ ������ � ������ �� ������. ����������������   � � ��������� ���������� ��������������� �������. ������� ��    ����� ������� ������!�r/P /Just L /Text ������ ��� �������  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0�    0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  �    ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  , �   rial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�1 �   1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�;  , A�     , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !��   ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,�   0 ,  0 , None , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 �   0 ,  0 ,  , !�;  , Arial ,  10 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �    0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 ,  0 ,  �     0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,  0 , �   ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�1  ,  ,  0 ,  0 ,  0 ,  0 ,�    ����������� ���������� ��������� � �������������� ������� �   � "List of all guests", � ��������� ��� ������� �� ������ (�    "Bills list for selected guest"). ���� � ����� "List of al�   l guests" ������ �����, �� � "Bills list for selected guest�   " ��������� ������ ���� ��� � ������ ��� ������. � ���������   � ������ ��������� ������ �� ���������� � ������ ������ ����   �� ����� �����.!�'/P /Just L /Text ������ �������� (Bill) �   ������������� ��� ������ � ������� � �� �������. ����� �����   ���� (Lists) ��������� ������������� ��������������� �������   . ������ �������� (Time) ������������� ��� ��������� � �����   ������� ���������� �� ������ � �����. ������� ����������� -M    �������� ������ � ��������������� ������� ���������� �� ��  ����� ���������, ����������� �������� ����� � ��������� ����   ���� ��������� ���������� ������� � ���� ������� ������� ���   ��� �������� �� ����� �������� �� ������ �������� (Bill). ��   ������� � ��������� � ���� ���������������. ��� ������� �����   ����. ����� ����� "Bills list for selected guest" ������� �  ���� ������ ���������� "Post edit" (F12);!�: /B /Just L /Te  xt �������� �� ������ ������ � ��� �� �����;!�. /B /Just L 6   /Text ���������� ��������� �������;!�) /B /Just L /Text ���  �������� ������ �������������� ���:!�= /B /Just L /Text ���h   ����� �������� �����:!��/B /Just L /Text ����� ����� � ��   - ��� ��������, ��������� � ��������������� ����. ��������  ��� ������ ����� ����� Rooms used.��������� �������� ������  , �� ����� ������������� ���������� ���������� ��������� ��	   ����� ������ ���������� ����� ��������� ��� ������ �������
  ���� ������� ������ ���� ���������� ������ �������. ���� ��  �������� ��������� ������� �� �����. ��������� ������ �����  � ������� � �������� ���� ��� ���������� ����� � ���������   /Link f:\work\guana_~1\gr\micros~1\myproj~1\guana\help\img\  ierh.wmf /Just L /Text ������������� ������������ ������ ��  ������ (Bill) �������� ��, ��� ����� �� ��� ������� ����� �<   ���� � ��������.!�� /P /Just L /Text ���������� ����������!  ����������� ������� ������ �� �������� ������).!��/P /Jus  ������� ���������� � ������� ������ "Post edit" �� �������   ���������� ����� (��� ������ �� ������������� ��� ���������   � ���������� ���������� ��� �������� �� ������ ������ � ��  ���� Exit;!�/B /Just L /Text ���������� ��������� �������  � ��������;!�6 /B /Just L /Text ���������� ���������� �� ��  ����� ���������� ���������:!�? /B /Just L /Text F2 - ������   �������������� ����������� ������;!�5 /B /Just L /Text ENT  ER - ����� �������������� ������;!�l /B /Just L /Text ESC -   ������ �������������� ������ (��������������� �������� ���  ������� ���� ����� ������);!�4 /B /Just L /Text F12 - �����  ����� ��������� ������.!�� /P /Just L /Text �������� �����  �� ESC ��� �������������� ������������ ������ � �����������   ��� ����� ����������� ����������. ��� ������� ESC � ������   �������������� ��� �� ���������� ����������� ������ ������0  t L /Text ��� ������� ������ �� �������� ������ ������� �  �� ������ ����� ��������� � ������ �����, �� ������ �������@  ����������.!�G /P /Just L /Text ���������� ����� ������� ��#  � ������������� �� ������ ����� � ������������ � ��������� $  ���������� ������ �������, �� ����� ����������� ������ ����%  ������ � ����� ����� ������������������. ���� �� ��������� &   ����� ��������, ��� ��� ���������� ����� ������� ��� �����'  �� �������������, ����������� �������� �������� ����������.(  ������� ������ �� ������-���� ��������. ��������� ����� ���)  l edit".!��/P /Just L /Text �� ���� ������ ����������� ���*  ���� ��������� �������� ESC, ���� ������� ���������� "Cance+  ���, ��������� ������. ��������� ��������� ������ ���� ����,  ����� ����� ��������������� �� ����� �� ��������� ����� ���-   ��� ������� �� ������ �������� ��� ���������� ����������. .  ������. ���������� ����� � ������� �� ������ ������ � �����/  �������� �� ������ � ���������� ���������� ���� ������ �����"  nav.wmf /Macro /Play /Popup /Just C!�j /P /Just L /Text ���3  ��� ���� ��������� ������ ������ �������� ���� '*'. �������4   ������ ����� � ����� ������ ���� ������ �� ��������� �����5  ��� ���������� ����� ������.!�= /P /Just L /Text ����� ����6  � ���������� � ���� ������� �����:!�v /B /Just L /Text ����7  ������� �� ������� (��������� ��������� �� ���������� �����8   ���������� � ����� ������ �� ������);!�} /B /Just L /Text 9  �������������� ����������� ������ (������� ���������� �����:  ���� ������������ ����� ��������� ������ ������).!�� /P /Ju;  st L /Text � ������� ���������� �� ������ ������ ����������<  �� �� �������, ������������� ��������� � ��������� ����� ��=  ����. ������ �� ����� ������� �� ��������� ��������� ������>  �����, ������� ��� ��������� ������� ������.!�i /I /Jump /L1  ink f:\work\guana_~1\gr\micros~1\myproj~1\guana\help\img\dbO  �� � ��������� ������ ����� ���������� ������ '*' � �������?  ���������� ����� ���������:!�� /B /Just L /Text ������ ����:2  ��� ������ (����� ����).!�� /P /Just L /Text � ������ ����Q  ����� ����� � ������, ���� ��� ��������� ������ � ����� �� B  �� ������ ���� �� ������ ������� ����� ��������. �������� �C  � � ������� �������� "drag and drop" �������������� �������D  ����� ��������� � ����� ������������ ���������. ��� �������E  �� ����� �������������. ��������� ��������� ������������ � F  Just L /Text �� ����� ������ �������� ������ ����� ��� ����G  �� ���������� ������� � �����, ��� ��� ���� ������.!�~/P /H  � ������ �������� ������ ������). ������ �� ������ ������ �I  �� ��������� ����� ������ �������� ��� ����������� ��������J   ������ ������ ��� �������� ������ ������ � ������ ����� (�K  ������ ������� ������ ������.!�� /P /Just L /Text ���������L  ��������� � ����������� ������ ������ � ����������� ��� ���M  �� ������ ������;!�~ /B /Just L /Text �������� ������ "+" �N  ���� �������� ������ "Post edit" ���������� ���� ��������� A  ������� ����);!�B /B /Just L /Text ����������� ������ �����6`  ���������� ������ �����.!� /H /Just M /Text ������������!�a  ���������� ��� ������ �� ������ ������ ������� ���������� �    5   � Additional charges grid                           S  W   m�  �  . 	9       � Topic@IDH_TimeWnd	  � 200V  ���� ������� � ���� ����� ����� �������� ������ ��� ��������   �������� ���������� �����. ���� ������� �����������, �� ��x   !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !��  �� �������� ��������� �� ������� � ������� �� ���������. ��X  � �������� �������� ������ �� ������������ � �� ����������Y  � ������� F12 ��� ���������� ������. ��� ���� �������������Z  ������������ ������ ��� ���������� ����� ������ ����� �����[  � ���������. ���� �� ������ ������� � ������ ����� ����� ��\  � ������ ���������� ��������� ���������� � ������� ������ �]  �� ������� "+" ����������. ��� ������������ ���������� ����^   ���������� ������ ������ � ������ ����� ������� ����������_  d/P /Just L /Text ��� ���������� ����� ������� � ����� ���p  �����. �� ���������, ����� ��� ������� ������ "Refresh" ���q  ������������ DBNavigator ������������ �� ����� ����� � ����A   �� ��� ������ ��������� ��������� ����������. ��������� � �c  ��� �� ������ ����� � ����� List of all guests ��� ������� d  ��� ������������� ����� �� ������ �������� ����� ������� �b  ator, ����������� ��������� �������� ��� ��������. ������ �y  ���� Search ���������� � ������ ������� ������������ ������g  ��� List of all guests. ��� ����� ����� ��������������� ���j  j~1\guana\help\img\dbnav.bmp /Just L /Text ��������𑒑����=   �!�� /R /Link f:\work\guana_~1\gr\micros~1\myproj~1\guana\hl  O~     �  �� 	_   -�   !�u /P /Just L /Text ���������m   ���� ����� "Bills list for selected guest". ��������� ����    �� ������������� ������ � �����.  
w �  � 1005           &  �M�� 
� / 6 K     � Topic@IDH_Comments  �      1   � List of all guests                                �  ������� ��� ��� ��������� ������� ���������� ����������� ���  ��� ����������.��!�� /R /Link f:\work\guana_~1\gr\micros~1\�  ���� ������, � ����� ������� � ���� �����.!�/B /Just L /r  ��������.  ����� ������������ � ������ ������, ���� �� ����s  � ���������� ��� ������� ������ Close. ������ �������� �� �t  ��� ��������, �� ������ �������� ��� �������� � ������� ���u  ils of bill for: "Fname Lname"). ���� �� ����������� ������v  � ������� � ��������� �����, ����������� ������ ����� (Deta�    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !z   �� �����. ���� ����� ���� � ������, �� �� ������ ������� �e  �� �������. ��� ������������� ���������� ������� ��� ������i  ������������!�g /R /Link f:\work\guana_~1\gr\micros~1\mypro{  g\grid.bmp /Just L /Text ����� ��� ������� � �����쑒������|  R /Link f:\work\guana_~1\gr\micros~1\myproj~1\guana\help\im}   �������� ����� (� ������� ������ ������ ���������).��!�� /~  ����� ���� ����������. ����� ������� '#' ��������� ��������  myproj~1\guana\help\img\ttl.bmp /Just L /Text ��������� ����  Text ���� ����� � ������ ���, �� ���� ��� ��������. ��� ����  ��� ��������� ������ � �������� ������������. ���� ����� ���  ���������� ��� ���������, � ������� ����������� �����, �����  ������� ������ ����� ����� Additional charges ����������� ��   �� �������������� �������� ����� ����� Rooms used. ��� ����  es, ���� ������ �� ������ ����� ����� Payments, ���� �������  ��� ���� ������ �� ����������� ����� ����� Additional Charg�  xt ����������� ���������� ������� �� �����. ���� ���� ������  ��� ����� �������� �� ������� �� ������).!�/B /Just L /Te�  ����� (��������� ���������� �� ������������ �� �������� ����  ���� ������. ����� � ������ �� ����� ������������ ����� ����  d guest. ���������� ������������ �������� ������������ �����  ����, ���� �������� ���� ����� ����� Bills list for selecte�  ��� ������ (������ New Bill>>), ������ ������� ��������� ���  � �� ������ ������� � ���������� ������, �� ������� ��������  �� ����� ��������������� �����������. ����� ���������� �����  ��� ���� ������ ������ �� ������ ������ ����� ����� Recomm�  �� �� ������� �����. ����� ��������, ��� �������� �������� �  �������� ��� �������� ����� "UnPay". ��� ���� ������ �������  �� Deposit received � Balance Due. � ����������� �� ������ �  �������� ������ ��������� � �������� ����� � ����������� ���  �������� ��������, �� ������ ����������� ���������� � ���� �  � � ��������������� �����.!�^/B /Just L /Text ����� ���� ��  ������� Balance Due � Deposit received ����� ���������������  ��� ������������� ������������ ����������� �����. ������� ��  t"). ��� ���� � ������ editbox'��, ����������� ����� ������  ������� ������������� � ����� "Bills list for selected gues�  rol" ��������� � �����������, ����� ���� �������� ������� (�  �������������� ����� ��������������� ��, ��� ������ "Pay en�  �� �� ���������� � ������ �� ��������� � �������� �����. � �  ���� ����� ������� ������������� �����. ��� ���� �� ��������  ended bill �� ������ �������� (Lists). ������� ���������� �:�  ������ �� ������� ����� �� �������� �������� (����� ����� "�  rges, Payments, Rooms used, List of all rooms, List of all �  guest cat, List of all bill category, Recommended bill, Lis�  t of all guest bills). � ����� ������ ������� � ��������� ��  ������� ���� ����� ������� '#' ������������ �������� ������f  � ��������� �����. � ���� ������ � ��� ����� ������ DBNavig�  ������� �������� (r). ��� ������ �������������� ���� (o). ��   ���������� �������� ����������� ���������� � �������� � ���  ������ ��� ������ - �� �� �� ������ �������������. ��� �����  ���� ������������� ������. � ��������� ������ ������� ���� �  ���� � ���������� �������. ����� ������ ����� ��������� ���  L /Text �� ����� ������ ������������ ������� ��� �����������   ������� �� ������ �� ����� ����������� �����.!��/P /Just �  �������� ������. ����� ������� ��������� �������� ������ ���  ������ "Rooms used" �������� ������ ������������ �� ������ �  List of all rooms" ������ ��������). � ���������������� �� �  f all guests, Bills list for selected guest, Additional cha�   ����� ������������ � ��������� �������� ���� ���������� ���  ��� ������� '#'. ������������ ����� �������� � �������� ����  �� ����� ��������� ���������� (�������, PgUp, PgDown, Home,�   End).!�) /P /Just L /Text ����� ������ ���� �����:!�M /B /P  Just L /Text ����������� �������� � �������������� ������ (�    �D�� 
0 1 8 Q     � Topic@IDH_MainWindow  �  �    �  	  � 1011   �  ��?`     �  �� J�     � Gen�  eral concepts�� Y�     �  �� 	i�  c-�   !�6 /T N /Ju�  st M /Text ��������� ������� � �������� ������!� /H /Just �  M /Text ���������!��/P /Just L /Text ������ � ������� �����  ���������� ���� ������������� ������������, ���������������  � ���������� ��� �������, ��������� ����� �������� �������    � ����� �� ��������� ��� �����.  
� �                    �  � ���� ����������. ��������� �������� ����������, ����� ����  ���� �������������� ������ � ������, �������� ����� (List o�  �� ���� � ���� ����� ���������� ��������. �������� ���������  ���, �� ������������� �������� � ��� ��� ����� � �� ��������  �.!�� /B /Just L /Text Category - ��������� �����. ����� ���  ������� ���������, ������������ � ���������� ������, ����� o  R   �  �  . 	9       � Topic@IDH_BillWnd	  � 200    �� �����, ��� ������ "Post edit" ����������.  
� �       �  ��� ������� ������������� ����� ���� ������ F12, �� ������ �  ��� ��������� � ���� ������ ����� Additional Charges, �� ���   ������� ������������� ����. �������, ���� ��������, �� ����  ������� ����� ������ ������ ����� ���������� ������ � �� ���  ��� ��������, ��� ���� �� ������������� ������ �����, �� ���  ������ � ��������� �����. ���� ����� �� �����, �� � ��� ����  ��� ������� ������� ������, ������� �������� ����������� ���   ��� �������������.!��/R /Link f:\work\guana_~1\gr\micros~�  1\myproj~1\guana\help\img\cur_rec.wmf /Just L /Text ������ �  ����� ������� ������� ������� ����� �� ����� �� � �����. ��  ���� ������� ��������������. ���� �� ����������� ��� �����  ze <= 20 )!�* /B /Just L /Text State - ���� ( size = 2 )!�4�   <= size <= 50 )!�1 /B /Just L /Text City - ����� ( 1 <= si�  ( 1 <= size <= 30 )!�4 /B /Just L /Text Address - ����� ( 1�  ize <= 30 )!�? /B /Just L /Text Last Name  - ������� ����� �  (Lists)!�; /B /Just L /Text First Name - ��� ����� ( 1 <= s�  �������� ����� ����� List of all guest cat ������ �������� �  /Just M /Text ������ ���� ������!�/P /Just L /Text � �����   ������ ����� ����������� ���� ��� - ��� ������ ���������. �  ���� �� ��������� �����, �� �� ������ ����� ��� � ������� ��  ������. ������ ����� ����� �� ������� �������� � ��� �������  �. ������������ ����� ���������� ����� �������� �������. ���   ������ �������� ����������� - �� ����� ���� ���� ������ � R  ����������� ������� � ���������.��� ������� ����������� ����  �� � ������ ����� ����� ����� ��������. ��� ������� � ������  ������������ ������ �� �������� ����������.����� �������� ���   all guests grid�� U�     �  �� 	e	  k-�   !�% /T N �  yments /Link /Macro /Play /popup /Just L /Text Payments!�I �  /L /Jump IDH_RoomsUsed /Link /Macro /Play /popup /Just L /T�  ext Rooms used!�Q /L /Jump IDH_Calc /Link /Macro /Play /pop�  up /Just L /Text Caliculating parameters!�H /L /Jump IDH_En�  rol /Link /Macro /Play /popup /Just L /Text Pay enrolment!��  L /L /Jump IDH_Wizard /Link /Macro /Play /popup /Just L /Te�  xt Wizards''Wizards!�H /L /Jump IDH_Sorte /Link /Macro /Pla�  y /popup /Just L /Text Sorting order!�@ /L /Jump IDH_Lists �  /Link /Macro /Play /popup /Just L /Text Lists!�_ /L /Jump I�  DH_ListBills /Link /Macro /Play /popup /Just L /Text List o    f all guest's bills (time)  
{ �                         +  ��� ������������� �������� ��� ������� ����� �����.!�b /L /!  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  �    ���� 
' - 4 M     � Topic@IDH_Guests  �    �  �  	  � 1007   �  ��;\     �  �� F�     � List of:�   /popup /Just L /Text Additional charges!�F /L /Jump IDH_Pa�  �������� ��� ������ ��������� �� �����, �� �� ������ �������  � ����� ���������� ������� �� ������ ��������� ������ � ����  ������ ����. ��� ��� ����� ������������� �������������� � �U  ����� ( date >= 1 ������ 1990 ).!�Y/P /Just L /Text �������  ��� ������������ ����� ������. ����� ����, ������� ���������  , ��� ���� �� ������ ���������� ����� ������������ ����� � �  ����� "Bills list for selected guest", �� ��� �� ���������   ���� ���� � ������� F12 ��� ������ �������, �� ���������� �     ,  0 ,  0 ,  0 ,  0 ,  0 ,  , !�                          �  Rules_for_DBGris /Link /Macro /Play /popup /Just L /Text Ru�  les of grids uning!�N /L /Jump IDH_Guests /Link /Macro /Pla�  y /popup /Just L /Text List of all guests!�[ /L /Jump IDH_B   illsLst /Link /Macro /Play /popup /Just L /Text Bills list k   ��     �  ��9V     �  �� @n     � IDH_Dubl�� �  for selected guest!�M /L /Jump IDH_AddCh /Link /Macro /Play�  ��� ��������� ������ �� ���������. ���� �� ����� ������� ��  �� ��������� � ������ ������ ���������� �����.!�b /L /Jump  ������� ������������������ - ���������� ���������� ������ �  ������� ���������� ������������ ������ (�����). ������� ���  ������ ���������� ���������, �� �� ����� ���� ��������� ��   ���� ������ � ���� �������).!�� /B /Just L /Text Name - ���  ����� ��������� ������. ������������ ��� ������� ������ ���	  ��� ������ ���������� ������ �������� ���������, �������� �
  ������ ����� �������� ����� ����� "List of all bill categor  y" �������� Lists.!�C /B /Just L /Text Amount - �������� ��  ��� ���������� (amount >= 0 ).!�L/B /Just L /Text Date - �  ��� ����������. ��� �������������� ���������. ���� �� ��� �  � �������, �� ��������� ��� �� ������ ��������� �������� ��  ������ �����, �� ������� �� ���������� ��������� ������� ��  �������� �� �����. ���� �� ��������� ������� ������ � �����  �������� �����, �� �������� ������� ������ ������� �� ��� ���   IDH_Rules_for_DBGris /Link /Macro /Play /popup /Just L /TeO   /B /Just L /Text Post - �������� ������ ( post > 0 )!�� /By  /P /Just L /Text ���������� ������� � ���� ����� ����� ����  ������ ��� ��������� � ������ ������ ���������� �����.!�  ���� ���������� ������������������ - ���������� ����������   ���� �� ������� ���������� ������������ ������ (�����). ���  ������ ������� ���������� ���������, �� �� ����� ���� �����  ������� ���� ���� � ������� F12 ��� ������ �������, �� ����  �, �� ����� ������������ ����� ������. ����� ����, �������    ������� �������� ���������� �����. ���� ������� ����������  t ���������� ������� � ���� ����� ����� �������� ������ ���   - �������� ������� ( 1 <= size <= 64 ).!�Y/P /Just L /Tex  ���������� �����. �� �������� ���������, ��� ������� ������+  �� ������ ������ ��� ����� � ������ ����. ����� �� �������    ��������, ��� ���� �� ������ ���������� ����� ������������   ����� � ����� "Bills list for selected guest", �� ��� �� ��0  �� ������ � ���� �������).!�8 /B /Just L /Text Amount - ���1  /B /Just L /Text Name room - �������� �������. ������, ����"  e to - ���� ������������  ( Date to >= 1 ������ 1990 ).!�� #  ��� ( Date from >= 1 ������ 1990 ).!�K /B /Just L /Text Dat$  Guests <= 50 ).!�K /B /Just L /Text Date from - ���� ������%  of Guests - ����� ������, ���������� ������� ( 0 <= No. of &   �� ������ ������ � ���� �������).!�_ /B /Just L /Text No. '  �� ��������� ���� ��������� (F12, 'Post edit", ���� �������(  , ��� �������������� ����� ���������� ������ ����� ��������)  ���� � ������������ ��� ������ � ������ editbox'�. �������*  ������ � ���� ������, �� ����� �������� ����������� �������-    �  	  � 1013   �  ��>_     �  �� I~     � Room.  s used grid�� X�     �  �� 	h%	  �-�   !�- /T N /Just/   M /Text ����� ������������� ������!��/P /Just L /Text ���  �� �� �� ������������ ������ ������, ���������� ������ ��   �� ������� ( amount >= 0 ).!�D /B /Just L /Text Description�@  ��� ���������� ��� ������� ������ � ������ �����, �������� A  ���� ����� � ����� "Bills list for selected guest", �� ��� 2  ���� ��������, ��� ���� �� ������ ���������� ����� ��������3  ������, �� ����� ������������ ����� ������. ����� ����, ���4  � ��� ������� �������� ���������� �����. ���� ������� �����5   /Text ���������� ������� � ���� ����� ����� �������� �����6   Rooms rate = Nights * No. of Guests * Charge!�Y/P /Just L7  ��.  ��� ���������� ����. ��� ������ ������������� ������. 8  �����.!�� /B /Just L /Text Charge - �������� ����� �� �����9  ��������� �� ������ ������ � ����������� �� ���� �������� �:   ������ ������������� ������. ��� �������� ����������� ����;  s rate - ����� �� ������� � ����.  ��� ���������� ����. ���<  ����. Nights = Date to - Date from!�� /B /Just L /Text Room=  ��� �����. ��� ���������� ����. ��� ������ ������������� ��>  l rooms" �� �������� Lists.!�y /B /Just L /Text Nights - ��?  �������� ������. ��� ����� �������� ����� ����� "List of al:P  �� ��������� ���� ���� � ������� F12 ��� ������ �������, ��Q   /B N /Just L /Text Total = Subtotal + [Tax+Service] - Paym�  ���� � �������. ��� ��������� ������������� ������, �������C  L /Text ����� �������� ��������� �������� ���������� ��� ��F  !  m�� 
/ - 4 M     � Topic@IDH_Wizard  �    G  �  	  � 1016   �  ��;\     �  �� Fs     � WizardsH  �� U�     �  �� 	e  �-�   !�d /P /Just L /Text ����I  ��������� ��� ��������� ���������� ����� ������ � ������. �J  ������ 2 ����������:!�& /B /Just L /Text ��� ���������� ���N  ��;!�& /B /Just L /Text ��� ���������� �����.!�� /P /Just L     Bill>>).  
| �                                          K  ��������� � ���������� ������ ����� ��� ����� �� ����� (NewL  ��. ����������� ���������� ������ ��������� ������������� �M   /Text ����������� ���� ����������� �������� ���������� ����   /Just L /Text Deposit - ������� ( deposit >= 0 ). ���� �� c   ���������� ������� ���������� ���������, �� �� ����� ���� �  ents!�g /B N /Just L /Text Deposit received - �����, ������S  � �� ������������ ������ �������� ���������� ����� �������T  ��� �����. �� �������� ��������� ��� ������� �������� �����U  � ������ ��� ����� � ������ ����. ����� �� ������� ������ �V   ���� ������, �� ����� �������� ����������� ����������� � �W  ����������� ��� ������ � ������ editbox'�. �������, ��� ��X  ������������ ����� ���������� ������ ����� ���������� �����!  ���� ���� ��������� (F12, 'Post edit", ���� ������� �� ����Z  �  ���� 
+ 7 > W     � Topic@IDH_Rules_for_DBGris[    �    �  	  � 1014   �  ��Ef     �  �� P�     \  � Rules for using DBGrids�� _�     �  �� 	o�  -�  #D   !�) /T N /Just M /Text Rules for using DBGris!�/P /Just ^  order�� T�     �  �� 	d�   ^ -�   !�T /P /Just L /Text_   ��������� ����������  �������� ���������� ������� ��������    �� �����.  
� �                                              04                                                         :R  /Text ����� �������� (payments)!��/P /Just L /Text ����� �q  . ������� ���������� ������������������ - ���������� ������b  ��������� �� ������� ���������� ������������ ������ (�����)�  Play /popup /Just L /Text General concepts!�Z /L /Jump IDH_f  al charges grid�� T�     �  �� 	d�  @-�   !�# /T N /g  Just M /Text ����� ����������!��/P /Just L /Text ����� ��h   �� ������������ ������ ���������� ���������� ����� �������i  ��� �����. �� �������� ��������� ��� ������� �������� �����j  � ������ ��� ����� � ������ ����. ����� �� ������� ������ �k   ���� ������, �� ����� ���������� ����������� ����������� �l   ������������ ��� ������ � ������ editbox'�. �������, ��� m  �������������� ����� ���������� ������ ����� ���������� ���  ������ ���� ��������� (F12, 'Post edit", ���� ������� �� ��o    G��� 
� / 6 O     � Topic@IDH_Payments  �  p    �  	  � 1012   �  ��=^     �  �� H{     � Paymea  nts grid�� W�     �  �� 	g�  i-�   !�, /T N /Just M :�  ���� ������ ��� ��������� � ������ ������ ���������� ������  ����� ������ ��� ��������� � ������ ������ ���������� ����r  ). ������� ���������� ������������������ - ���������� �����s   ��������� �� ������� ���������� ������������ ������ (�����t  � ���������� ������� ���������� ���������, �� �� ����� ����u  � ��������� ����� ����� � ������� F12 ��� ������ �������, �v   ������������ ����� � ����� "List of all guestst", �� ��� �w  ���, ������� ��������, ��� ���� �� ������ ���������� ������x  ���� ������ ��� ������� �������� ���������� �����.  ����� �  ��� ����� � ������ ������ �������� ������� (�� ������������z  �/P /Just L /Text �� ������ ������� ���������, ��� ������ {    	 !�1 /T N /Just M /Text ������ ������ ���������� �����!�|   list for selected guest grid�� W�     �  �� 	g�  -�}    �  	  � 1002   �  ��=^     �  �� H�   '  �" Bills    p /Just L /Text ��. ������� ������ � �������  
� �         .!�b /L /Jump IDH_Rules_for_DBGris /Link /Macro /Play /popu�/  �.!�b /L /Jump IDH_Rules_for_DBGris /Link /Macro /Play /pop�  ���������� ������ ����� ���������� �������� ���� ����������   �������� F12 ��� ������ ��������.!�F /B N /Just L /Text To�  tal additional = Sum( Additional Charges.Amount )!�: /B N /�  Just L /Text Total payments = Sum( Payments.Amount )!�= /B �  N /Just L /Text Total rooms = Sum( Rooms Used.Rooms rate )!�  �< /B N /Just L /Text Subtotal = Total additional + Total rB  ooms!�0 /B N /Just L /Text Tax+Service = 17% �� Subtotal!�>�   � �������� ����� ��� ���������� ������� (Pay enrol)!�� /B �  N /Just L /Text Balance Due - �����, ������� ����� ������� �  ������ ����� �������� � ��� ���������. ���� �� �������� ���    �� �� �������, �� ��� ����� > 0, ����� 0.  
� �          �  � Balance Due ����������.!��/B /Just L /Text �������� �����  ��������� ������� ����� Deposit received �� ������� �����, �  �   �b�� 
 , 3 L     � Topic@IDH_Sorte  �    �]    	  � 1015   �  ��:[     �  �� Ex     � Sorting :�  ayments", "Rooms used". �������, ��� ���������� ���� ����� �  ������� � �������� � ��������� � Deposit received, � �������  �� Total - Deposit received ��������� � Balance Due. ��� ���  ������ ����������� ������ ����������.!�� /B /Just L /Text ��  ������ ����� � ������ ���������� �� ����� (������ UnPay). ��  ������������� ��������� ������� �������� ����� ���� �������  ����/��������� �����. ������ ��������� ����� ������ ��������  ���� �� ������� �����. ��� ����� �� ������ ������� ������� �  ������ Deposit ����� "List of all guests" (������� ����) � �  /P /Just L /Text �� ������ ������ �������� ����������� �����  �������� ��� ������. ���� ������ ������.!�) /B /Just L /Te�  T  	�� 
� + 2 K     � Topic@IDH_Calc  �    � �   	  � 1003   �  ��9Z     �  �� D�   $  � Calculati�  ng parameters of Bills�� S�     �  �� 	cK  �-�  	 !��  /P N /Just L /Text ������������� ����������� �� ������, ���  ����� ��� �������� ����� � ������ "Additional Charges", "P6�  ��� �� �������� Total � �������� ��� ��������. ��� ����� ���   L /Text ��������� ������;!�T /B /Just L /Text �������� ����   �������;!�" /B /Just L /Text ��������� ������;!�" /B /Just�  �!�" /P /Just L /Text ������� 4 ������:!� /B /Just L /Text�  ���� ������ �� ������ �� �������� �� ������, ������� ��� ���  ���������, �� ���������� ���������� �������;!�j /B /Just L �  �� ����������� ��� ��������� ������������ �����.!�8/P /Jus�  ��� ������ "UnPay", �� ������ - "Pay enrol". ���������� ����  ������ ��� �� ����������� ���������. � ������ ������ �������  t L /Text ����� ��������, ��� ���� ������ ��������� � ������  ����� �������� ���������� ��� ������ � ��������.!�� /P /Jus�  ���� �������� ������, ����������� ������ ����� ����� � �����  ������ ����� ���������-�������� ������� �� ����������. ��� �  �������� 3 ��������:!�o/B /Just L /Text ���������� ������ �  ����� �� ����� (�������� ������ Pay enrol). ��� ���� �������  ����� �����, ������� ����� ���� ����� � �������� �����, ���6�  ������ ��������� ������ ��� ������ �� ��������� ������.!�d �  �������� ������� ��������� ������, �� ������� ��������������  � ����������� ������ � ��������� ��������� ���������. ����     ��. ������� ������ � �������  
� �                       �  ��������� ������������� ��� ���� ���������� ������ ���������  �  ���� 
. , 3 L     � Topic@IDH_Enrol  �    ��    +�� 
, , 3 L     � Topic@IDH_Lists  �    ��    	  � 1009   �  ��:[     �  �� Ep   
  � Lists���   T�     �  �� 	d  �-�   !� /T N /Just M /Text ������  ������ �������� ���������. ���� ������ ��������� ������.!�)�  Text �� ������ ��������� ������ �������� ����������� �������  ) /B /Just L /Text Name ( 1 <= size <= 30 )!� /P /Just L /�  ������� �������� ���������. ���� ������ ��������� ������.!��  /Text �� ������ ��������� ������ �������� ����������� ������  �� �� ������� � ���� ( 0 <= Rate <= 100000 )!� /P /Just L �  xt Name ( 1 <= size <= 40 )!�H /B /Just L /Text Rate - ����    xt ��. ������� ������ � �������  
� �                    �   ���������� ������ �� ���������� ��������� � ��������� �����   ������� ��, ��� � ������ ������ ������������ � �����. ����  �������������� �������� ������ "Remove all". ��� ���� ������  ������ ����������� ��� �������� ���������� ������ �� ����. �  �����������.!�~/P /Just L /Text ��������� �������� ������ �  �� Bill � ���������� ������������� ����� � ������������ ����   ������ ������ <<Jump to, ��� ������� � �������� �� �������  ���". ��� �������������� �� ������ ������� � ����� ������ ��  �.!�� /P /Just L /Text ����� ��������� � ������ "������ ����  �������� �������� ������ �� ���� �� ��������� ���� ���������  ���� ��� ��������� ��������� ������;!�P /B /Just L /Text ���  /Text ���������� �� ���� ������ �� ��������� ���������� ����   /Just L /Text ������������ ���:!�~ /B /Just L /Text �������   !�0 /T N /Just M /Text ��������������� ������ ������!�" /P�   of all guest's bills grid�� X�     �  �� 	h*  �-�  �  �� ����������� ���������������� �������� ���������� �� �����  ����� "Refill" ��� ���������� ������ ���������.!�/P /Just�  ��� "Lists", �� ����� �������� �� �������� "Time" ������� ��  xt ���� �� ��������������� ������ ��������� ������ �� ������  ��������� � ��������� � ������ ���������.!�� /P /Just L /Te�  ���� ����� ������������ ����� ������ ��� ������, ������� ���   � ������������ ����� ������ ���� ���������. � ��������� ���  �����-������ "All guests" ��������, �� ���� ������ ���������  /Just M /Text ������ ��������� ������!�b/P /Just L /Text ��  goryes filtering�� X�     �  �� 	h  i-�   !�* /T N �    �  	  � 1010   �  ��>_     �  �� I�     � Cate�    ���� 
 0 7 P     � Topic@IDH_LstFltCat  �  �    ?O�� 
� + 2 G     � Topic@IDH_Dubl  �    �     ooments button                                            �  H_Rules_for_DBGris /Link /Macro /Play /popup /Just L /Text �   �� �������� (From, To � ������� ���������).!�b /L /Jump ID�   L /Text ����� ��������, ��� ������ "Print" (������ � ������   � �� �������� ��������� ���������. ����� �������� ����� ���   ������ "Rooms used" ������� ����� ������������ ����� ����,�  �����  ���� ����, �� ���  ��� ��������� ����� ����������� ��  ������ ����� ����� �������� ������ �� ������������ � �� ���  y enrol". ������, ������� �������, ��� ����  �� �����  �����  ��������� "UnPay", �������� �������� ������ � ��������� "Pa�  ������, Additional Charges) ��� ��� ������������ �����, �� �  t L /Text ���� �� ������ �������� �������� ������ ����� (���    	  � 1006   �  ��:[     �  �� E{     � Making e�  nrolment�� T�     �  �� 	d�  Z-�   !�3 /T N /Just M �  /Text �������� �� ������� � ����������!�% /P /Just L /Text     guests" ������ ������ ���������.  
� �                   �  � �������� �� ����������. ��� ���������� ������������ "All �  ������� ��������� ������ ��� ��� ������ ������ �������������  ��� ������) ��������� ������ � ������ ���� ���� ������� ���   � ����� ���������� � ������ "Rooms used" ����� �� ������� �  ������� � �������� � � ���� ������, ������������� �� � ����  ��� ���� ���������. ���� �� ������ �������� ���������, �� ��  �� ���� ����� ���� ���������. ������� �� ������ ������� ����  , �� �� ������ ������� ��������� ������, ���� � ������ �����  ����� ������ ������� ������������ � ������ ������. ���������  ��� �� �� ������ ������� �������, ��������� ������ ��� �����  me ( 1 <= size <= 30 )!��/P /Just L /Text ����� ��������, �  ext ���� ������ ������������� �����.!�) /B /Just L /Text Na�   /B /Just L /Text Name ( 1 <= size <= 25 )!�1 /P /Just L /T&  	  ��� 
� , 3 L     � Topic@IDH_Enrol  �    �    ������� ������ � "List of Rooms" �������� "Lists".  
� � �  ��� � ��������� "Pay enrol". ����� ������������ �������� ��  ������ ��������� ���� �������� ��������� ������ ����� ������  "List of Rooms" �������� "Lists". ����� ����� �� ������ ����   ���� "Rooms rate" � ������ � � ������ ������ ����� ����� :  ��� ������. ���������� ��� ��������� �������.!�� /P /Just L  (date >= 1 ������ 1990).!�M /B /Just L /Text Folio - �����   ��� ������.!�D /B /Just L /Text Date - ���� �������� �����   ������� ����� ����� ���� ������ ������, ������� � ����� ���  Bill no - ����� �����. �������� ���������� ���������������   �������� ��������� ������ ���� ������.!�� /B /Just L /Text   ���� ����������� ������������ ������ �����. ��������������   �� ������" ��� ������� ������ ������� �����. �� ������ ����  �������� � ���� textbox'�� � ������ �������� � ������ "����	  ��� ���� ������ ������ ������� ��� �����. ���� ����� ������
  �� ����� ����� �� ������ ���� �������, ��� ������������ ���   � ����� � ��������� �����, ����������� ������ �����). ����.  ���.!�b /L /Jump IDH_Rules_for_DBGris /Link /Macro /Play /p  � ��� ����������� ������� ������������ ������ ��������� ���  ���� �� �������. ���� �� � ��������, �� ��� �� ��������� �   /Text ���������� �� ������� ���������� �������� �������� �   ����� ������������� ����� ( 1 <= size <= 15 ).!�3 /B /Just     Gris>!�  !�  !�  !�  !�                                      H_Rules_for_DBGris>!�) ������,(Global), 0,<IDH_Rules_for_DB  (Global), 2,<IDH_Rules_for_DBGris>!�( �����,(Global), 2,<ID    �  ��     �  ��=Z     �  �� Dv     � IDH_Comme  nts�� S�     �  �� 	c  � -�   !�x /P /Just L /Text �  �������� ������������� ����� ����������� � ���������� �����`  . ���� ����������� �������� ��������������.  
 �  � 10�  F   Td  � ) 	0       � Topic@Topic1  �    � C    ust L /Text ��. ������� ������ � �������  
� �              /L /Jump IDH_Rules_for_DBGris /Link /Macro /Play /popup /J  ������� ����� � ������� textbox'���), � �� ����� �����.!�b  ������� � �������� ����� ������ Comments (��������� ����� �  ents - ( 1 <= size <=256 ). ��� ���� �� ����������� ��� ���  ext Details - ( 1 <= size <= 64 ).!�� /B /Just L /Text Comm  L /Text Heard of GI - ( 1 <= size <= 35 ).!�/ /B /Just L /T    !�  !�  !�  !�  !�  !�  !�  !�  !�  !�                                                                                    "                                                             #                                                             $                                                             %                                                             (  �  .0�� 
( , 3 L     � Topic@IDH_AddCh  �    �e    	  � 1001   �  ��:[     �  �� E�     � Addition~  �  %��� 
* / 6 O     � Topic@IDH_BillsLst  �       /Text ��. ������� ������ � �������  
� �                *  Jump IDH_Rules_for_DBGris /Link /Macro /Play /popup /Just L-  3  o��� 
- 0 7 P     � Topic@IDH_ListBills  �  �    �  	  � 1008   �  ��>_     �  �� I�   #  � List    opup /Just L /Text ��. ������� ������ � �������  
y �        up /Just L /Text ��. ������� ������ � �������  
� �      ,  .	  ���� 
) 0 7 P     � Topic@IDH_RoomsUsed  �  